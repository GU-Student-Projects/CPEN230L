<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-53.5564,10.9668,89.3936,-63.2832</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-35.5,-14.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-35.5,-18.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-35.5,-22</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>-16.5,-14.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>-16.5,-19.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>-16.5,-24.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND3</type>
<position>3,-7.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND3</type>
<position>3,-16</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>15 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_NAND3</type>
<position>3,-23.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>12 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>-22,-13.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>-22,-18.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>-22,-23.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>-30.5,-14.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>-30.5,-18.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>-30.5,-22</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>31</ID>
<type>DE_TO</type>
<position>-11,-14.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>32</ID>
<type>DE_TO</type>
<position>-11,-19.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>33</ID>
<type>DE_TO</type>
<position>-11,-24.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>-2.5,-5.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>-2.5,-16</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>-2.5,-25.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>-2.5,-7.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>-2.5,-9.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>-2.5,-18</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>-2.5,-14</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>-2.5,-21.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>-2.5,-23.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>44</ID>
<type>BA_NAND4</type>
<position>17.5,-15.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>24 </input>
<input>
<ID>IN_3</ID>27 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>23.5,-15.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>BA_NAND4</type>
<position>3,-32</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>IN_3</ID>29 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>-4,-29</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>-4,-33</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>-4,-35</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-2,0</position>
<gparam>LABEL_TEXT Gabe DiMartino, September 18, 2023</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,-13.5,-19.5,-13.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-19.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-19.5,-15.5,-19.5,-13.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,-23.5,-19.5,-23.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-19.5,-25.5,-19.5,-23.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,-18.5,-19.5,-18.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-19.5,-20.5,-19.5,-18.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33.5,-14.5,-32.5,-14.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33.5,-18.5,-32.5,-18.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33.5,-22,-32.5,-22</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-14.5,-13,-14.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-19.5,-13,-19.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-24.5,-13,-24.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-5.5,0,-5.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-16,0,-16</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-25.5,0,-25.5</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-7.5,0,-7.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>0 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>0,-7.5,0,-7.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-9.5,0,-9.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>0 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>0,-9.5,0,-9.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-18,0,-18</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-0.5,-14,0,-14</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>0 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>0,-14,0,-14</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-21.5,0,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-23.5,0,-23.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-12.5,10,-7.5</points>
<intersection>-12.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-12.5,14.5,-12.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-7.5,10,-7.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-16,10,-14.5</points>
<intersection>-16 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-14.5,14.5,-14.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-16,10,-16</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-15.5,22.5,-15.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-23.5,10,-16.5</points>
<intersection>-23.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-16.5,14.5,-16.5</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-23.5,10,-23.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-29,0,-29</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-2 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-2,-31,-2,-29</points>
<intersection>-31 4</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-2,-31,0,-31</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-2 2</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-32,11.5,-18.5</points>
<intersection>-32 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-32,11.5,-32</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-18.5,14.5,-18.5</points>
<connection>
<GID>44</GID>
<name>IN_3</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2,-33,0,-33</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2,-35,0,-35</points>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,190.6,-99</PageViewport></page 1>
<page 2>
<PageViewport>0,0,190.6,-99</PageViewport></page 2>
<page 3>
<PageViewport>0,0,190.6,-99</PageViewport></page 3>
<page 4>
<PageViewport>0,0,190.6,-99</PageViewport></page 4>
<page 5>
<PageViewport>0,0,190.6,-99</PageViewport></page 5>
<page 6>
<PageViewport>0,0,190.6,-99</PageViewport></page 6>
<page 7>
<PageViewport>0,0,190.6,-99</PageViewport></page 7>
<page 8>
<PageViewport>0,0,190.6,-99</PageViewport></page 8>
<page 9>
<PageViewport>0,0,190.6,-99</PageViewport></page 9></circuit>