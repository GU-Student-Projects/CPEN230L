<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-24.3064,10.9668,118.644,-63.2832</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>10.5,-24.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>10.5,-27.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>15,-24.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>15,-27.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>38,-26</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>32,-25</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>32,-27</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>42,-26</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>56.5,-25</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>56.5,-27</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>66.5,-26</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR2</type>
<position>62,-26</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>73,-26</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_INVERTER</type>
<position>78.5,-26</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>83,-26</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>BA_NAND2</type>
<position>29.5,-36.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>BA_NAND2</type>
<position>37,-36.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>24,-35.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>24,-37.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>42,-36.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>BA_NAND2</type>
<position>54,-33.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>BA_NAND2</type>
<position>54,-39</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>BA_NAND2</type>
<position>61.5,-36.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>48.5,-33.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>48.5,-39</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>66.5,-36.5</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>BA_NAND2</type>
<position>78,-36.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>72.5,-36.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>83,-36.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>BE_NOR2</type>
<position>54,-46.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>BE_NOR2</type>
<position>61.5,-46.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>66.5,-46.5</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>48.5,-45.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>48.5,-47.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>23.5,-43.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>23.5,-49</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>41.5,-46</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>BE_NOR2</type>
<position>29.5,-43.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>BE_NOR2</type>
<position>29.5,-49</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>BE_NOR2</type>
<position>36,-46</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>72.5,-46.5</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>66</ID>
<type>BE_NOR2</type>
<position>78,-46.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>83,-46.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>13,-34.5</position>
<gparam>LABEL_TEXT NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>13,-45</position>
<gparam>LABEL_TEXT NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>13,-37.5</position>
<gparam>LABEL_TEXT Implementation</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>12.5,-48</position>
<gparam>LABEL_TEXT Implementation</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>40,-19.5</position>
<gparam>LABEL_TEXT A*B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>64.5,-19.5</position>
<gparam>LABEL_TEXT A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>82.5,-20</position>
<gparam>LABEL_TEXT A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>45,-13</position>
<gparam>LABEL_TEXT Gabe DiMartino, September 18, 2023</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-24.5,13,-24.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>13 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>13,-24.5,13,-24.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-27.5,13,-27.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>34,-25,35,-25</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>34,-27,35,-27</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-26,41,-26</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-26,41,-26</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>65,-26,65.5,-26</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>58.5,-25,59,-25</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>58.5,-27,59,-27</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>75,-26,75.5,-26</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>81.5,-26,82,-26</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-36.5,34,-36.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>34 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>34,-37.5,34,-35.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-35.5,26.5,-35.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>26,-37.5,26.5,-37.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>40,-36.5,41,-36.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>37</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>51,-34.5,51,-32.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-33.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-33.5,51,-33.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>51 2</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>51,-40,51,-38</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-39 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-39,51,-39</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>51 2</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-35.5,57.5,-33.5</points>
<intersection>-35.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-35.5,58.5,-35.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-33.5,57.5,-33.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-39,57.5,-37.5</points>
<intersection>-39 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-37.5,58.5,-37.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-39,57.5,-39</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-36.5,65.5,-36.5</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>41</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>75,-37.5,75,-35.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-36.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>74.5,-36.5,75,-36.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-36.5,82,-36.5</points>
<connection>
<GID>47</GID>
<name>N_in0</name></connection>
<connection>
<GID>45</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-47.5,58.5,-45.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-46.5,58.5,-46.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-46.5,65.5,-46.5</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-45.5,51,-45.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-47.5,51,-47.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-45,32.5,-43.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-45,33,-45</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-49,32.5,-47</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-47,33,-47</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-46,40.5,-46</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-44.5,26,-42.5</points>
<intersection>-44.5 3</intersection>
<intersection>-43.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-42.5,26.5,-42.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-43.5,26,-43.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-44.5,26.5,-44.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-50,26,-48</points>
<intersection>-50 3</intersection>
<intersection>-49 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-49,26,-49</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-48,26.5,-48</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-50,26.5,-50</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-47.5,74.5,-45.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-47.5 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-45.5,75,-45.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-47.5,75,-47.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-46.5,82,-46.5</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<connection>
<GID>66</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,190.6,-99</PageViewport></page 1>
<page 2>
<PageViewport>0,0,190.6,-99</PageViewport></page 2>
<page 3>
<PageViewport>0,0,190.6,-99</PageViewport></page 3>
<page 4>
<PageViewport>0,0,190.6,-99</PageViewport></page 4>
<page 5>
<PageViewport>0,0,190.6,-99</PageViewport></page 5>
<page 6>
<PageViewport>0,0,190.6,-99</PageViewport></page 6>
<page 7>
<PageViewport>0,0,190.6,-99</PageViewport></page 7>
<page 8>
<PageViewport>0,0,190.6,-99</PageViewport></page 8>
<page 9>
<PageViewport>0,0,190.6,-99</PageViewport></page 9></circuit>