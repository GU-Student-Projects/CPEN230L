<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-53.5564,10.9668,89.3936,-63.2832</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-25,-8.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-25,-14.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-25,-20</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>-5,-8.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>-5,-14.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>-5,-20.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND3</type>
<position>10,-14.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>18.5,-14.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>-20.5,-8.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>-20.5,-14.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>-20.5,-20</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>-12.5,-7.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>-12.5,-13.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>-12.5,-9.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>-12.5,-15.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>-12.5,-21.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>-12.5,-19.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-25,-6</position>
<gparam>LABEL_TEXT SW1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-25,-12</position>
<gparam>LABEL_TEXT SW2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>-25,-18</position>
<gparam>LABEL_TEXT SW3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>-9.5,-6</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>-9.5,-8.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>-9.5,-12.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>-9.5,-14.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>-9.5,-18</position>
<gparam>LABEL_TEXT 9</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>-0.5,-9.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>-0.5,-15.5</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>-9.5,-20.5</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>-0.5,-21.5</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>5.5,-11.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>5.5,-13.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>5.5,-15.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>15,-15.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>0,-7.5</position>
<gparam>LABEL_TEXT U1A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>0,-13.5</position>
<gparam>LABEL_TEXT U1B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>0,-19.5</position>
<gparam>LABEL_TEXT U1C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>15,-13.5</position>
<gparam>LABEL_TEXT U2A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>-3.5,-25.5</position>
<gparam>LABEL_TEXT U1: 7400 Quad 2-input NAND, VCC pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>-3.5,-27.5</position>
<gparam>LABEL_TEXT U2: 7410 Triple 3-input NAND, VCC pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>-3,-30</position>
<gparam>LABEL_TEXT Switches and LEDs correspond to Logic Trainer I/O devices</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>-4,-2.5</position>
<gparam>LABEL_TEXT Gabe DiMartino, September 18, 2023</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>-3.5,1</position>
<gparam>LABEL_TEXT H = ((AB)'*(AC)'*(BC)')'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>21.5,-14</position>
<gparam>LABEL_TEXT H</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-12.5,2,-8.5</points>
<intersection>-12.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-12.5,7,-12.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-8.5,2,-8.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-14.5,7,-14.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-20.5,2,-16.5</points>
<intersection>-20.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-16.5,7,-16.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-20.5,2,-20.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-14.5,17.5,-14.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,-8.5,-22.5,-8.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,-14.5,-22.5,-14.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22.5,-14.5,-22.5,-14.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,-20,-22.5,-20</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-7.5,-8,-7.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-13.5,-8,-13.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-9.5,-8,-9.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-15.5,-8,-15.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-21.5,-8,-21.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-19.5,-8,-19.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,190.6,-99</PageViewport></page 1>
<page 2>
<PageViewport>0,0,190.6,-99</PageViewport></page 2>
<page 3>
<PageViewport>0,0,190.6,-99</PageViewport></page 3>
<page 4>
<PageViewport>0,0,190.6,-99</PageViewport></page 4>
<page 5>
<PageViewport>0,0,190.6,-99</PageViewport></page 5>
<page 6>
<PageViewport>0,0,190.6,-99</PageViewport></page 6>
<page 7>
<PageViewport>0,0,190.6,-99</PageViewport></page 7>
<page 8>
<PageViewport>0,0,190.6,-99</PageViewport></page 8>
<page 9>
<PageViewport>0,0,190.6,-99</PageViewport></page 9></circuit>