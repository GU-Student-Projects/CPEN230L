<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-3.62216,0.439692,82.7918,-48.7236</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>46.5,-34.5</position>
<gparam>LABEL_TEXT chosen Y input</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>33.5,-21.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>9 </output>
<input>
<ID>SEL_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>13,-25</position>
<gparam>LABEL_TEXT 0 or 1 for X, 0 to 3 for Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_MUX_4x1</type>
<position>34.5,-34.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>11 </input>
<output>
<ID>OUT</ID>8 </output>
<input>
<ID>SEL_0</ID>1 </input>
<input>
<ID>SEL_1</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>29,-20.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>29,-22.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>29,-37.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>29,-33.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>29,-35.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>29,-31.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>39,-34.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>39,-21.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>DD_KEYPAD_HEX</type>
<position>18.5,-16</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>2 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>17,-23</position>
<gparam>LABEL_TEXT MUX address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>26.5,-20.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>26.5,-22.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>26.5,-31.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>26.5,-33.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>26.5,-37.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>26.5,-35.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>35,-17</position>
<gparam>LABEL_TEXT 1-bit wide 2-to-1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>35,-27</position>
<gparam>LABEL_TEXT 1-bit wide 4-to-1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>34,-7</position>
<gparam>LABEL_TEXT A MUX chooses between inputs.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>49,-38</position>
<gparam>LABEL_TEXT (See pages 2-4 for more.)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>46,-21.5</position>
<gparam>LABEL_TEXT chosen X input</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-28.5,23.5,-19</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-28.5 2</intersection>
<intersection>-19 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-28.5,35.5,-28.5</points>
<intersection>23.5 0</intersection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-29.5,35.5,-28.5</points>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23.5,-19,33.5,-19</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-29.5,24.5,-17</points>
<intersection>-29.5 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-17,24.5,-17</points>
<connection>
<GID>20</GID>
<name>OUT_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-29.5,34.5,-29.5</points>
<connection>
<GID>4</GID>
<name>SEL_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-20.5,31.5,-20.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-22.5,31.5,-22.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>31,-33.5,31.5,-33.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>12</ID>
<points>31,-37.5,31.5,-37.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>37.5,-34.5,38,-34.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-21.5,38,-21.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>17</ID>
<points>31,-31.5,31.5,-31.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>31,-35.5,31.5,-35.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>15.0882,-11.3632,101.503,-60.5268</PageViewport>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>51.5,-50.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>27.5,-45.5</position>
<gparam>LABEL_TEXT 0 to 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>81,-41.5</position>
<gparam>LABEL_TEXT chosen Y input</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>58.5,-23</position>
<gparam>LABEL_TEXT from gates</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>51.5,-37.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>51.5,-44</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>51.5,-31</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>39</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-36.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<output>
<ID>OUT_1</ID>15 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>28,-44</position>
<gparam>LABEL_TEXT MUX Address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>49,-31</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>49,-37.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>49,-50.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>49,-44</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AE_SMALL_INVERTER</type>
<position>38,-40</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_SMALL_INVERTER</type>
<position>38,-44.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>42.5,-40</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1'</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>42.5,-37.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>42.5,-44.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0'</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>42.5,-42</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>58.5,-27</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>58.5,-29</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>58.5,-33.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>58.5,-35.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0'</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>58.5,-40</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1'</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>58.5,-42</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>58.5,-46.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1'</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>58.5,-48.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0'</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND3</type>
<position>64,-29</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>33 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND3</type>
<position>64,-35.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<input>
<ID>IN_2</ID>34 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND3</type>
<position>64,-42</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<input>
<ID>IN_2</ID>35 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND3</type>
<position>64,-48.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>36 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR4</type>
<position>71,-39</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>76.5,-39</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>59.5,-20.5</position>
<gparam>LABEL_TEXT 1-bit wide 4-to-1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-50.5,61,-50.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-42,40.5,-42</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>34 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>34,-44.5,34,-39.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 23</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>34,-44.5,36,-44.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>34 7</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-37.5,40.5,-37.5</points>
<connection>
<GID>39</GID>
<name>OUT_1</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>35 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35,-40,35,-37.5</points>
<intersection>-40 12</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>35,-40,36,-40</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>35 5</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>22</ID>
<points>40,-40,40.5,-40</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>40,-44.5,40.5,-44.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-27,61,-27</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-29,61,-29</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-35.5,61,-35.5</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-33.5,61,-33.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-40,61,-40</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-42,61,-42</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>60.5,-46.5,61,-46.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-31,61,-31</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-37.5,61,-37.5</points>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-44,61,-44</points>
<connection>
<GID>88</GID>
<name>IN_2</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>60.5,-48.5,61,-48.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-36,68,-29</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-29,68,-29</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-38,67,-35.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-38,68,-38</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-42,67,-40</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-40,68,-40</points>
<connection>
<GID>91</GID>
<name>IN_2</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-48.5,68,-42</points>
<connection>
<GID>91</GID>
<name>IN_3</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67,-48.5,68,-48.5</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-39,75.5,-39</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<connection>
<GID>93</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>16.7391,-4.28689,108.838,-56.6843</PageViewport>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>50,-40.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>67.5,-14</position>
<gparam>LABEL_TEXT 1-bit wide 4-to-1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>50,-31.5</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>50,-36</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>50,-27</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>97</ID>
<type>DD_KEYPAD_HEX</type>
<position>40,-20.5</position>
<output>
<ID>OUT_0</ID>64 </output>
<output>
<ID>OUT_1</ID>65 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>29,-20.5</position>
<gparam>LABEL_TEXT Address (0 to 3)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>47.5,-27</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>47.5,-31.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>47.5,-40.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>47.5,-36</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AE_OR4</type>
<position>68,-34.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>77 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>123</ID>
<type>GA_LED</type>
<position>73.5,-34.5</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>BA_DECODER_2x4</type>
<position>50.5,-22</position>
<input>
<ID>ENABLE</ID>66 </input>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT_0</ID>67 </output>
<output>
<ID>OUT_1</ID>68 </output>
<output>
<ID>OUT_2</ID>69 </output>
<output>
<ID>OUT_3</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>EE_VDD</type>
<position>46.5,-19.5</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>61,-28</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND2</type>
<position>61,-32.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_AND2</type>
<position>61,-37</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_AND2</type>
<position>61,-41.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>67.5,-17</position>
<gparam>LABEL_TEXT from a 2-to-4 decoder and gates</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>42.5,-33</position>
<gparam>LABEL_TEXT Inputs</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>78,-36.5</position>
<gparam>LABEL_TEXT chosen Y input</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-40.5,58,-40.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-34.5,72.5,-34.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-23.5,47.5,-23.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>45,-21.5,47.5,-21.5</points>
<connection>
<GID>97</GID>
<name>OUT_1</name></connection>
<intersection>47.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>47.5,-22.5,47.5,-21.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-21.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-20.5,47.5,-20.5</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-42.5,54,-23.5</points>
<intersection>-42.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-42.5,58,-42.5</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-23.5,54,-23.5</points>
<connection>
<GID>125</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-38,55,-22.5</points>
<intersection>-38 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-22.5,55,-22.5</points>
<connection>
<GID>125</GID>
<name>OUT_1</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-38,58,-38</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-33.5,56,-21.5</points>
<intersection>-33.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-21.5,56,-21.5</points>
<connection>
<GID>125</GID>
<name>OUT_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-33.5,58,-33.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-29,57,-20.5</points>
<intersection>-29 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-20.5,57,-20.5</points>
<connection>
<GID>125</GID>
<name>OUT_3</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-29,58,-29</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-27,58,-27</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-31.5,58,-31.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-36,58,-36</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-41.5,65,-37.5</points>
<connection>
<GID>122</GID>
<name>IN_3</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64,-41.5,65,-41.5</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-37,64,-35.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-35.5,65,-35.5</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-33.5,64,-32.5</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-33.5,65,-33.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-31.5,65,-28</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64,-28,65,-28</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-3.60739,-5.65694,82.8061,-54.82</PageViewport>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>49.5,-20.5</position>
<gparam>LABEL_TEXT from 4 1-bit wide 2-to-1 MUXs</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_MUX_2x1</type>
<position>36,-31</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>82 </output>
<input>
<ID>SEL_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_MUX_2x1</type>
<position>36,-37</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>81 </output>
<input>
<ID>SEL_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_MUX_2x1</type>
<position>36,-43</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>80 </output>
<input>
<ID>SEL_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_MUX_2x1</type>
<position>36,-49</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>79 </output>
<input>
<ID>SEL_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>DD_KEYPAD_HEX</type>
<position>19,-14.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<output>
<ID>OUT_1</ID>89 </output>
<output>
<ID>OUT_2</ID>90 </output>
<output>
<ID>OUT_3</ID>91 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>165</ID>
<type>DD_KEYPAD_HEX</type>
<position>19,-27</position>
<output>
<ID>OUT_0</ID>84 </output>
<output>
<ID>OUT_1</ID>85 </output>
<output>
<ID>OUT_2</ID>86 </output>
<output>
<ID>OUT_3</ID>87 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>167</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>43,-40.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>81 </input>
<input>
<ID>IN_3</ID>82 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_TOGGLE</type>
<position>18.5,-46.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>11,-46</position>
<gparam>LABEL_TEXT Address (0 or 1)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>11,-14.5</position>
<gparam>LABEL_TEXT Input 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>11,-26</position>
<gparam>LABEL_TEXT Input 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>50.5,-17.5</position>
<gparam>LABEL_TEXT 4-bit wide 2-to-1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-49,39.5,-41.5</points>
<intersection>-49 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-41.5,40,-41.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-49,39.5,-49</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-43,38.5,-40.5</points>
<intersection>-43 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-40.5,40,-40.5</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-43,38.5,-43</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-39.5,38.5,-37</points>
<intersection>-39.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-39.5,40,-39.5</points>
<connection>
<GID>167</GID>
<name>IN_2</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-37,38.5,-37</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-38.5,39.5,-31</points>
<intersection>-38.5 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-38.5,40,-38.5</points>
<connection>
<GID>167</GID>
<name>IN_3</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-31,39.5,-31</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-46.5,32.5,-28.5</points>
<intersection>-46.5 1</intersection>
<intersection>-40.5 57</intersection>
<intersection>-34.5 56</intersection>
<intersection>-28.5 55</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-46.5,36,-46.5</points>
<connection>
<GID>161</GID>
<name>SEL_0</name></connection>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>32.5,-28.5,36,-28.5</points>
<connection>
<GID>155</GID>
<name>SEL_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>32.5,-34.5,36,-34.5</points>
<connection>
<GID>157</GID>
<name>SEL_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>32.5,-40.5,36,-40.5</points>
<connection>
<GID>159</GID>
<name>SEL_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-50,24.5,-30</points>
<intersection>-50 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-50,34,-50</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-30,24.5,-30</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-44,34,-44</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>25 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>25,-44,25,-28</points>
<intersection>-44 1</intersection>
<intersection>-28 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>24,-28,25,-28</points>
<connection>
<GID>165</GID>
<name>OUT_1</name></connection>
<intersection>25 6</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-38,25.5,-26</points>
<intersection>-38 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-38,34,-38</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-26,25.5,-26</points>
<connection>
<GID>165</GID>
<name>OUT_2</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-32,26,-24</points>
<intersection>-32 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-32,34,-32</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-24,26,-24</points>
<connection>
<GID>165</GID>
<name>OUT_3</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-48,28.5,-17.5</points>
<intersection>-48 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-48,34,-48</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-17.5,28.5,-17.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-42,29,-15.5</points>
<intersection>-42 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-42,34,-42</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-15.5,29,-15.5</points>
<connection>
<GID>163</GID>
<name>OUT_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-36,29.5,-13.5</points>
<intersection>-36 3</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-13.5,29.5,-13.5</points>
<connection>
<GID>163</GID>
<name>OUT_2</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-36,34,-36</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-30,30,-11.5</points>
<intersection>-30 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-30,34,-30</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-11.5,30,-11.5</points>
<connection>
<GID>163</GID>
<name>OUT_3</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-20.5906,92.7576,626.783,-275.551</PageViewport></page 4>
<page 5>
<PageViewport>-55.6686,144.26,807.494,-346.817</PageViewport></page 5>
<page 6>
<PageViewport>-55.6686,144.26,807.494,-346.817</PageViewport></page 6>
<page 7>
<PageViewport>-55.6686,144.26,807.494,-346.817</PageViewport></page 7>
<page 8>
<PageViewport>-55.6686,144.26,807.494,-346.817</PageViewport></page 8>
<page 9>
<PageViewport>-55.6686,144.26,807.494,-346.817</PageViewport></page 9></circuit>