<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-64.4608,5.9178,208.944,-134.014</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>31,-63</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_OR2</type>
<position>31.5,-76</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>31.5,-91</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>32,-26.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>BE_NOR2</type>
<position>31.5,-40.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_INVERTER</type>
<position>31,-53</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>43,-63</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>43,-76</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>43,-91</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>43.5,-26.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>43.5,-40.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>43.5,-53</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>46.5,-26</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>47,-40</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>47,-52.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>47,-62.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>46.5,-75.5</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>46,-90.5</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>8.5,-55</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>8.5,-60</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>9,-50</position>
<gparam>LABEL_TEXT SW1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>8.5,-64</position>
<gparam>LABEL_TEXT SW2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>26.5,-23</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>26,-37</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>26,-50</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>26,-59.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>26,-72.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>26,-87.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>26.5,-29</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>26,-43.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>26,-66</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>26,-78.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>26,-94.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>36,-28.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>36,-43</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>36.5,-54.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>35,-65</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>35.5,-77.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>35,-93</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>38,-24.5</position>
<gparam>LABEL_TEXT U1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>37.5,-38.5</position>
<gparam>LABEL_TEXT U2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>37.5,-50.5</position>
<gparam>LABEL_TEXT U3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>36.5,-60.5</position>
<gparam>LABEL_TEXT U4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>37,-74</position>
<gparam>LABEL_TEXT U5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>37,-89</position>
<gparam>LABEL_TEXT U6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>86,-31.5</position>
<gparam>LABEL_TEXT U1: 7400	Quad 2-input NAND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>85,-46.5</position>
<gparam>LABEL_TEXT U2: 7402	Quad 2-input NOR, Vcc pin 14, Gnd pin 7</gparam>
<gparam>Quad 2-input NAND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>83,-58</position>
<gparam>LABEL_TEXT U3: 7404 Hex Inverters, Vcc pin 14, Gnd pin 7 </gparam>
<gparam>Quad 2-input NAND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>87,-70</position>
<gparam>LABEL_TEXT U4: 7408 Quad 2-input AND, Vcc pin 14, Gnd pin 7 </gparam>
<gparam>Quad 2-input NAND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>86,-83.5</position>
<gparam>LABEL_TEXT U5: 7432 Quad 2-input OR, Vcc pin 14, Gnd pin 7 </gparam>
<gparam>Quad 2-input NAND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>87.5,-96</position>
<gparam>LABEL_TEXT U6: 7486 Quad 2-input XOR, Vcc pin 14, Gnd pin 7 </gparam>
<gparam>Quad 2-input NAND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>54,-107.5</position>
<gparam>LABEL_TEXT Switches and LEDs correspond to Logic Trainer I/O devices</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>57.5,-17.5</position>
<gparam>LABEL_TEXT Gabe DiMartino, September 11, 2023</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>24,-6.5</position>
<gparam>LABEL_TEXT A = (SW1*SW2)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>24.5,-12</position>
<gparam>LABEL_TEXT B = (SW1+SW2)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>46.5,-6.5</position>
<gparam>LABEL_TEXT C = SW1'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>50,-12</position>
<gparam>LABEL_TEXT D = SW1*SW2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>73,-6.5</position>
<gparam>LABEL_TEXT E = SW1+SW2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>86,-12</position>
<gparam>LABEL_TEXT F = (SW1*SW2') + (SW1'*SW2) </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-63,42,-63</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-76,42,-76</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-91,42,-91</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-26.5,42.5,-26.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-40.5,42.5,-40.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>22</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-53,42.5,-53</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-55,19.5,-25.5</points>
<intersection>-55 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-25.5,29,-25.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection>
<intersection>22 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-55,19.5,-55</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22,-90,22,-25.5</points>
<intersection>-90 5</intersection>
<intersection>-75 6</intersection>
<intersection>-62 7</intersection>
<intersection>-53 8</intersection>
<intersection>-39.5 9</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>22,-90,28.5,-90</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>22 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>22,-75,28.5,-75</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>22 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22,-62,28,-62</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>22 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>22,-53,28,-53</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>22 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22,-39.5,28.5,-39.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>22 4</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-92,19.5,-60</points>
<intersection>-92 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-60,19.5,-60</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-92,28.5,-92</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection>
<intersection>23.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-92,23.5,-27.5</points>
<intersection>-92 2</intersection>
<intersection>-77 9</intersection>
<intersection>-64 8</intersection>
<intersection>-41.5 7</intersection>
<intersection>-27.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>23.5,-27.5,29,-27.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>23.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>23.5,-41.5,28.5,-41.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>23.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>23.5,-64,28,-64</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>23.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>23.5,-77,28.5,-77</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>23.5 3</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 1>
<page 2>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 2>
<page 3>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 3>
<page 4>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 4>
<page 5>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 5>
<page 6>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 6>
<page 7>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 7>
<page 8>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 8>
<page 9>
<PageViewport>0,238.236,1778,-671.764</PageViewport></page 9></circuit>