<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-8.94734,24.5614,48.3114,-47.0121</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>21,-13</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>18,-6</position>
<gparam>LABEL_TEXT E = SW1*SW2 + SW3*SW4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>24.5,-11</position>
<gparam>LABEL_TEXT U1A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>35,-14</position>
<gparam>LABEL_TEXT U2A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>21.5,-27</position>
<gparam>LABEL_TEXT U1: 7408 Quad 2-Input AND, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>21,-22</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>21,-29</position>
<gparam>LABEL_TEXT U2: 7432 Quad 2-Input OR, Vcc pin 14, Gnd pin 7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>17.5,-10.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>40,-17.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>17.5,-15</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>24.5,-14</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>32,-17.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>17.5,-19</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>17.5,-24</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>42.5,-17</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>24.5,-23</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>7,-11</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>19,-8</position>
<gparam>LABEL_TEXT Gabe DiMartino, September 5, 2023</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>7,-15</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>7,-20</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>28.5,-13</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>7,-23.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>29,-21.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>29,-15</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>3.5,-11</position>
<gparam>LABEL_TEXT SW1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>29,-19.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>4,-14.5</position>
<gparam>LABEL_TEXT SW2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>35,-16.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>4,-19.5</position>
<gparam>LABEL_TEXT SW3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>31,-12.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>4,-23.5</position>
<gparam>LABEL_TEXT SW4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>31.5,-21.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>24.5,-20.5</position>
<gparam>LABEL_TEXT U1B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>22.5,-32</position>
<gparam>LABEL_TEXT Switches and LEDs correspond to Logic Trainer I/O devices.</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-12,13.5,-11</points>
<intersection>-12 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-12,18,-12</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-11,13.5,-11</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-15,13.5,-14</points>
<intersection>-15 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-14,18,-14</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-15,13.5,-15</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-21,13.5,-20</points>
<intersection>-21 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-20,13.5,-20</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-21,18,-21</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-23.5,18,-23.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>18 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-23.5,18,-23</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-16.5,26.5,-13</points>
<intersection>-16.5 1</intersection>
<intersection>-13 2</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-16.5,29,-16.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-13,27.5,-13</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-22,26.5,-18.5</points>
<intersection>-22 2</intersection>
<intersection>-21.5 3</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-18.5,29,-18.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-22,26.5,-22</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-21.5,28,-21.5</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-17.5,39,-17.5</points>
<connection>
<GID>15</GID>
<name>N_in0</name></connection>
<connection>
<GID>19</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 1>
<page 2>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 2>
<page 3>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 3>
<page 4>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 4>
<page 5>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 5>
<page 6>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 6>
<page 7>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 7>
<page 8>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 8>
<page 9>
<PageViewport>0,374.799,696,-495.201</PageViewport></page 9></circuit>